library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity hex2sseg is
    Port ( hex : in STD_LOGIC_VECTOR (3 downto 0);
           sseg : out STD_LOGIC_VECTOR (6 downto 0));
end hex2sseg;

architecture Behavioral of hex2sseg is

begin


end Behavioral;
